-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 17.1.0 Build 590 10/25/2017 SJ Lite Edition
-- Created on Sat Dec 23 14:29:31 2017

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY loadSignalGen IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        CS : OUT STD_LOGIC;
        Din : OUT STD_LOGIC;
        freezeParalell : OUT STD_LOGIC
    );
END loadSignalGen;

ARCHITECTURE BEHAVIOR OF loadSignalGen IS
    TYPE type_fstate IS (Origin,state1,state2,state3,state4,state5,state6,state7,state8,state9,state10,state11,state12,state13,state14,state15,state16,state17,state18,state20,state21,state23,state22,state24,state19);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= Origin;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate)
    BEGIN
        CS <= '0';
        Din <= '0';
        freezeParalell <= '0';
        CASE fstate IS
            WHEN Origin =>
                reg_fstate <= state1;

                Din <= '0';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state1 =>
                reg_fstate <= state2;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state2 =>
                reg_fstate <= state3;

                Din <= '0';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state3 =>
                reg_fstate <= state4;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state4 =>
                reg_fstate <= state5;

                Din <= '0';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state5 =>
                reg_fstate <= state6;

                Din <= '0';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state6 =>
                reg_fstate <= state7;

                Din <= '0';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state7 =>
                reg_fstate <= state8;

                Din <= '0';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state8 =>
                reg_fstate <= state9;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state9 =>
                reg_fstate <= state10;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state10 =>
                reg_fstate <= state11;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state11 =>
                reg_fstate <= state12;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state12 =>
                reg_fstate <= state13;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state13 =>
                reg_fstate <= state14;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state14 =>
                reg_fstate <= state15;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state15 =>
                reg_fstate <= state16;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state16 =>
                reg_fstate <= state17;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state17 =>
                reg_fstate <= state18;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state18 =>
                reg_fstate <= state19;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state20 =>
                reg_fstate <= state21;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state21 =>
                reg_fstate <= state22;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state23 =>
                reg_fstate <= state24;

                Din <= '1';

                freezeParalell <= '1';

                CS <= '0';
            WHEN state22 =>
                reg_fstate <= state23;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN state24 =>
                reg_fstate <= state24;

                Din <= '1';

                freezeParalell <= '1';

                CS <= '1';
            WHEN state19 =>
                reg_fstate <= state20;

                Din <= '1';

                freezeParalell <= '0';

                CS <= '0';
            WHEN OTHERS => 
                CS <= 'X';
                Din <= 'X';
                freezeParalell <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
