--Write comparator function.