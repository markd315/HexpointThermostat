/*Write comparator function.